module mmu(

);


endmodule